../struct_from_matlab/tb.sv