../dpi_c_ex_types.svh