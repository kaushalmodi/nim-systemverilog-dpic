../dpi_c_ex_test.sv