// Time-stamp: <2019-02-26 12:48:37 kmodi>

program top;

  import "DPI-C" hello=task hello();

  initial begin
    hello();
  end

endprogram : top
