// Time-stamp: <2019-01-17 21:59:34 kmodi>

program top;

  import "DPI-C" hello=task hello();

  initial begin
    hello();
  end

endprogram
