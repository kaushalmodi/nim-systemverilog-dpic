../svvpi/sv/vpi_pkg.sv