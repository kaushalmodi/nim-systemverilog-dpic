orig/test.sv