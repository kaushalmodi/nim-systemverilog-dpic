orig/amiq_top.sv