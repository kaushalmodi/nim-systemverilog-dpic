../tb.sv