// Time-stamp: <2014-11-17 23:27:09 kmodi>

// Source: http://www.testbench.in/DP_03_IMPORT.html

program main;

   import "DPI-C" string_sv2c=task string_sv2c();

      initial begin
         string_sv2c();
      end

endprogram
